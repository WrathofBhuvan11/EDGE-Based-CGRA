// g_tile.sv
// Global control tile: Manages block fetching, commitment, speculation (up to 8 in-flight blocks), branch handling with EXIT_ID, morph configuration propagation (e.g., revitalization for S-morph), and debug signals.
// Instantiates block_controller for atomicity and termination detection (constant outputs via header mask).
// Hierarchy: Standalone with block_controller sub-module; interfaces to external control_if and internal instr_fetch_if.
// G-tile fetches block addr to I-tile, tracks in-flight, speculation/multiblock;
//     - Commit/dealloc on completion/flush; Revitalization signal for S-morph loops, 
//     - Block execution flow, constant outputs/store mask for termination;
//     - Branches with EXIT_ID for multiple exits

`include "includes/trips_defines.svh"
`include "includes/trips_types.svh"
`include "includes/trips_interfaces.svh"
`include "includes/trips_isa.svh"
`include "includes/trips_params.svh"
`include "includes/trips_config.svh"

module g_tile (
    input clk,                                    // Clock input
    input rst_n,                                  // Reset input (active-low)
    input morph_config_t morph_config,            // Morph configuration input (D/T/S modes)
    // External control_if ports (master: outputs fetch/commit signals)
    output logic fetch_req,                       // Fetch request output to external (part of control_if.master)
    output logic [31:0] block_addr,               // Block address output for fetch 
    input logic commit,                           // Block commit input signal
    input logic branch_taken,                     // Branch outcome input
    output logic [(`MAX_INFLIGHT_BLOCKS-1):0] block_id,  // In-flight block ID output (up to 8)
    output logic revitalize,                      // Revitalization output for S-morph loops
    // Internal instr_fetch_if ports (master: to I-tile for fetch)
    output logic instr_fetch_req,                 // Internal fetch request to I-tile 
    output logic [31:0] instr_block_addr,         // Internal block address to I-tile
    input instr_t [(`BLOCK_SIZE-1):0] instructions,  // Instructions input from I-tile (up to 128)
    input block_header_t header,                  // Block header input (store mask etc)
    input logic ready,                            // Fetch ready input from I-tile
    // Debug outputs
    output logic debug_commit,                    // Debug commit output
    output logic [31:0] debug_pc                  // Debug current PC output
);

    // Internal signals
    logic [(`MAX_INFLIGHT_BLOCKS-1):0] inflight_blocks;  // Bitmap for in-flight blocks (speculation tracking)
    logic speculation_flush;                             // Flush signal on mispredict/mis-exit
    logic [4:0] exit_id_internal;                        // Internal EXIT_ID from branch 

    // Morph-specific logic (e.g., revitalize only in S-morph)
    assign revitalize = (morph_config.revitalize_enable) && (morph_config.morph_mode == `MORPH_S) && commit;  // Trigger on commit in S-morph

    // Assign external control_if outputs (master mode)
    assign block_addr = next_block_addr;                                   // Output predicted addr
    assign block_id = inflight_blocks;                                      // Output active IDs

    // Assign internal internal instr_fetch_if outputs (master to I-tile)
    assign instr_fetch_req = fetch_req;                                    // Mirror external fetch
    assign instr_block_addr = block_addr;                                  // Mirror addr

    // Debug: Commit from input, PC from current block_addr
    assign debug_commit = commit;
    assign debug_pc = block_addr;

    logic [31:0] next_block_addr;        // Next predicted block addr(for fetch)

    // Instantiate block_controller (for atomicity, termination, speculation flush)
    block_controller block_controller_inst (
        .clk(clk),
        .rst_n(rst_n),
        .morph_config(morph_config),                // Pass morph for frame/revitalization mgmt
        .commit(commit),                            // Input commit signal
        .branch_taken(branch_taken),                // Input branch outcome
        .exit_id(exit_id_internal),                 // Input EXIT_ID from branch instr
        .header(header),                            // Input block header (store mask/reg writes)
        .fetch_req(fetch_req),                      // Output fetch_req (generated by FSM)
        .ready(ready),                              // Input ready from I-tile
        .block_addr(block_addr),                    // Pass internal instr_block_addr as current base
        .inflight_blocks(inflight_blocks),          // Output in-flight bitmap
        .speculation_flush(speculation_flush),      // Output flush on mispredict
        .next_block_addr(next_block_addr)           // Output next predicted addr
    );

    // Speculation logic: Track in-flight, flush on mispredict (simplified FSM)
    typedef enum logic [1:0] {IDLE, FETCHING, EXECUTING, COMMITTING} state_t;
    state_t state, next_state;

    always_ff @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            state <= IDLE;
            inflight_blocks <= 0;
            exit_id_internal <= 0;  // Reset
        end else begin
            state <= next_state;
            if (fetch_req) inflight_blocks <= {inflight_blocks[`MAX_INFLIGHT_BLOCKS-2:0], 1'b1};  // Shift in new block
            if (commit) inflight_blocks <= inflight_blocks >> 1;  // Commit oldest
            if (speculation_flush) inflight_blocks <= inflight_blocks & 1'b1;  // Flush all but oldest
        end
    end

    always_comb begin
        next_state = state;
        case (state)
            IDLE: if (fetch_req) next_state = FETCHING;
            FETCHING: if (ready) next_state = EXECUTING;
            EXECUTING: if (commit) next_state = COMMITTING;
            COMMITTING: next_state = IDLE;
        endcase
        if (speculation_flush) next_state = IDLE;  // Override on flush
    end

    // Need to check - Branch/EXIT_ID handling: Update next_addr on taken (simplified; assume from branch instr via internal sig)
    // Need to check - Revitalization: Already assigned; broadcast to res stations via morph_config (in e_tile)
endmodule
